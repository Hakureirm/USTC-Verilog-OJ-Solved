module top_module(
    input a, 
    input b,
    output out );

    and a1(out,a,b);
endmodule
