module top_module( 
    input a, 
    input b, 
    output out );

    nor a1(out,a,b);
endmodule