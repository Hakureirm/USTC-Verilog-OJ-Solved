module top_module(
    input in, output out
);
    wire in,out;
    assign out = in;
endmodule